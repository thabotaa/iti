module AHMED  #(parameter ahmed#=2 