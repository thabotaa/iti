module AHMED_tb(); parameter ahmed#=2 